library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;    -- Biblioteca IEEE para funções aritméticas

entity ULA is
    generic
    (
        larguraDados : natural := 8
    );
    port
    (
      entradaA, entradaB:  in STD_LOGIC_VECTOR((larguraDados-1) downto 0);
      seletor:  in STD_LOGIC_VECTOR(2 downto 0);
      saida:    out STD_LOGIC_VECTOR((larguraDados-1) downto 0);
		flagLess : out std_logic;
      flagZero: out std_logic
    );
end entity;

architecture comportamento of ULA is
  --constant zero : std_logic_vector(larguraDados-1 downto 0) := (others => '0');

   signal soma :      STD_LOGIC_VECTOR((larguraDados-1) downto 0);
   signal subtracao : STD_LOGIC_VECTOR((larguraDados-1) downto 0);
   signal op_and :    STD_LOGIC_VECTOR((larguraDados-1) downto 0);
   signal op_or :     STD_LOGIC_VECTOR((larguraDados-1) downto 0);
   signal op_xor :    STD_LOGIC_VECTOR((larguraDados-1) downto 0);
   signal op_not :    STD_LOGIC_VECTOR((larguraDados-1) downto 0);
	
	signal A_extended : STD_LOGIC_VECTOR(larguraDados downto 0);
	signal B_extended : STD_LOGIC_VECTOR(larguraDados downto 0);
	signal subtracao_extended : STD_LOGIC_VECTOR(larguraDados downto 0);

    begin
		
		A_extended(larguraDados) <= '0';
		A_extended((larguraDados-1) downto 0) <= entradaA;
		
		B_extended(larguraDados) <= '0';
		B_extended((larguraDados-1) downto 0) <= entradaB;
	 
	 
      soma      <= STD_LOGIC_VECTOR(unsigned(entradaA) + unsigned(entradaB));
      subtracao <= STD_LOGIC_VECTOR(unsigned(entradaA) - unsigned(entradaB));
      op_and    <= entradaA and entradaB;
      op_or     <= entradaA or entradaB;
      op_xor    <= entradaA xor entradaB;
      op_not    <= not entradaA;
		subtracao_extended <= STD_LOGIC_VECTOR(signed(A_extended) - signed(B_extended));

      saida <= soma when (seletor = "000") else
          subtracao when (seletor = "001") else
          entradaA when  (seletor = "010") else
          entradaB when  (seletor = "011") else
          op_xor when    (seletor = "100") else
          op_not when    (seletor = "101") else
          op_and when    (seletor = "110") else
          op_or when     (seletor = "111") else
          entradaA;      -- outra opcao: saida = entradaA

      --flagZero <= '1' when unsigned(saida) = unsigned(zero) else '0';
      flagZero <= '1' when unsigned(saida) = 0 else '0';
		flagLess <= '1' when subtracao_extended(larguraDados) = '1' else '0';

end architecture;